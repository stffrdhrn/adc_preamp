* Components used to implement/simulate the ports for
* the preamp schematic. 

.INCLUDE UA741.301
*               + - G O V
.SUBCKT uA741CP 1 2 3 4 5
*      + - V G O
  XUI1 1 2 5 3 4 UA741
.ENDS uA741CP

* simulates a microphone at 10mV 440hz
.SUBCKT MIC_IN 1 2 3
  Vmic  1 3 ac SIN(0 0.02 440)
.ENDS MIC_IN

.SUBCKT OUT 1 2
  Rload 1 2 2K
.ENDS OUT

.SUBCKT PWR 1 2 3
  V1 2 1 DC 3.3v
  V2 3 1 DC 12v
.ENDS PWR

* D1n5819 from http://www.onsemi.com/pub_link/Collateral/1N5819.LIB
.MODEL DIODESCH D 
+IS=1.19279e-05 RS=0.0625421 N=1.16517 EG=1.3
+XTI=3.22098 BV=40 IBV=0.001 CJO=1.50114e-10
+VJ=1.5 M=0.590203 FC=0.5 TT=2.6273e-08
+KF=0 AF=1
