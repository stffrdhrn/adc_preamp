* EESchema Netlist Version 1.1 (Spice format) creation date: Wed 04 Feb 2015 22:25:01 JST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

.include components.cir

XU1  1 6 0 9 2 uA741CP		
R5  6 7 50K		
C1  4 1 4.7uF		
R6  9 7 1K1		
C3  9 8 10nF		
R7  8 0 18K		
R4  6 3 1K1		
C2  3 0 4.7uF		
R2  2 1 56K		
R3  1 0 56K		
R1  2 4 56K		
XJ1  0 0 4 JACK_2P		

*.op
*.ac dec 10 1 1e10
*.plot ac vdb(1), vdb(8)

.tran 0.1m 5m
.plot tran v(1), v(8)

.end
