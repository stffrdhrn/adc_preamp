* EESchema Netlist Version 1.1 (Spice format) creation date: Wed 06 May 2015 09:59:38 AM JST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0
.include components.cir

*Sheet Name:/
XU1  10 9 0 8 5 uA741CP		
R5  9 7 50K		
C1  2 10 4.7uF		
R6  8 7 1K1		
R7  1 0 18K		
R4  9 6 1K1		
C2  6 0 4.7uF		
R2  5 10 56K		
R3  10 0 56K		
R1  5 2 56K		
XJ1  2 0 0 MIC_IN		
C3  8 1 4.7uF		
R8  3 1 18K		
D2  1 3 DIODESCH		
D1  0 1 DIODESCH		
XP1  0 1 OUT		
XP2  0 3 5 PWR		

*.op
*.ac dec 10 1 50K
*.plot ac vdb(1), vdb(8)

.tran 0.1ms 5ms
.plot tran v(2), V(8), V(1)

.end
